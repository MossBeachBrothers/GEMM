//Top module for GEMM
module GEMM #()(

);


endmodule 


