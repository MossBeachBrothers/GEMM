//GEMM Controller Module

module GEMMController #()(

);

endmodule


