module SRAM #(parameter ADDR_WIDTH = 16, DATA_WIDTH =32)(

);

endmodule 

